//-----------------------------------------------------------------------------
// Project name: Verification of APB Protocol
// Version: 1.0
// Description: Package file for APB Protocol
// Author: Mehul Prajapati
//-----------------------------------------------------------------------------

package apb_pkg;

	`include "apb_trans.sv"
	`include "apb_gen.sv"
	`include "apb_drv.sv"
	`include "apb_mon.sv"
	`include "apb_sco.sv"
	`include "apb_env.sv"

endpackage