`ifndef AFIFO_DEFINES_SV
`define AFIFO_DEFINES_SV

`define WIDTH 8
`define DEPTH 16

`endif