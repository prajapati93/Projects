////////////////////////////////////////////////
// RAM Verification in SV
// File description: Defines RAM Size
// Author Name: Mehul Prajapati
// Version: 1.0
/////////////////////////////////////////////////

`ifndef RAM_DEFINES_SV
`define RAM_DEFINES_SV

`define ADDR_WIDTH 4
`define DATA_WIDTH 8

`endif