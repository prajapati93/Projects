////////////////////////////////////////////////
// FIFO Verification in SV
// File description: Package file
// Author Name: Mehul Prajapati
// Version: 1.0
/////////////////////////////////////////////////

package fifo_pkg;

	`include "fifo_trans.sv"
	`include "fifo_gen.sv"
	`include "fifo_driver.sv"
	`include "fifo_monitor.sv"
	`include "fifo_rf.sv"
	`include "fifo_sb.sv"
	`include "fifo_env.sv"

endpackage